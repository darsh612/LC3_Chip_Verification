//----------------------------------------------------------------------
// Created with uvmf_gen version 2022.3
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// DESCRIPTION: This class records data_mem transaction information using
//       a covergroup named data_mem_transaction_cg.  An instance of this
//       coverage component is instantiated in the uvmf_parameterized_agent
//       if the has_coverage flag is set.
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
class data_mem_transaction_coverage  extends uvm_subscriber #(.T(data_mem_transaction ));

  `uvm_component_utils( data_mem_transaction_coverage )

  T coverage_trans;

  // pragma uvmf custom class_item_additional begin
  // pragma uvmf custom class_item_additional end
  
  // ****************************************************************************
  covergroup dmem_txn_cg;
    // pragma uvmf custom covergroup begin
    // UVMF_CHANGE_ME : Add coverage bins, crosses, exclusions, etc. according to coverage needs.
    option.auto_bin_max=1024;
    option.per_instance=1;
    // complete_data: coverpoint coverage_trans.complete_data;
    // Data_dout: coverpoint coverage_trans.Data_dout;
    // Data_din: coverpoint coverage_trans.Data_din;
    // Data_rd: coverpoint coverage_trans.Data_rd;
    // Data_addr: coverpoint coverage_trans.Data_addr;
    Data_din: coverpoint coverage_trans.Data_din{
      bins _data = {[1:$]};
    }
    Data_rd: coverpoint coverage_trans.Data_rd
    {
    }
    Data_dout: coverpoint coverage_trans.Data_dout{
      bins  _data_dout = {0};
    }
    complete_data: coverpoint coverage_trans.complete_data;
    // pragma uvmf custom covergroup end
  endgroup

  // ****************************************************************************
  // FUNCTION : new()
  // This function is the standard SystemVerilog constructor.
  //
  function new(string name="", uvm_component parent=null);
    super.new(name,parent);
    dmem_txn_cg=new;
    // `uvm_warning("COVERAGE_MODEL_REVIEW", "A covergroup has been constructed which may need review because of either generation or re-generation with merging.  Please note that transaction variables added as a result of re-generation and merging are not automatically added to the covergroup.  Remove this warning after the covergroup has been reviewed.")
  endfunction

  // ****************************************************************************
  // FUNCTION : build_phase()
  // This function is the standard UVM build_phase.
  //
  function void build_phase(uvm_phase phase);
    dmem_txn_cg.set_inst_name($sformatf("dmem_txn_cg%s",get_full_name()));
  endfunction

  // ****************************************************************************
  // FUNCTION: write (T t)
  // This function is automatically executed when a transaction arrives on the
  // analysis_export.  It copies values from the variables in the transaction 
  // to local variables used to collect functional coverage.  
  //
  virtual function void write (T t);
    `uvm_info("COV","Received transaction",UVM_HIGH);
    coverage_trans = t;
    dmem_txn_cg.sample();
  endfunction

endclass

// pragma uvmf custom external begin
// pragma uvmf custom external end


// //----------------------------------------------------------------------
// // Created with uvmf_gen version 2022.3
// //----------------------------------------------------------------------
// // pragma uvmf custom header begin
// // pragma uvmf custom header end
// //----------------------------------------------------------------------
// //----------------------------------------------------------------------
// //     
// // DESCRIPTION: This class records data_mem transaction information using
// //       a covergroup named data_mem_transaction_cg.  An instance of this
// //       coverage component is instantiated in the uvmf_parameterized_agent
// //       if the has_coverage flag is set.
// //
// //----------------------------------------------------------------------
// //----------------------------------------------------------------------
// //
// class data_mem_transaction_coverage  extends uvm_subscriber #(.T(data_mem_transaction ));

//   `uvm_component_utils( data_mem_transaction_coverage )

//   T coverage_trans;

//   // pragma uvmf custom class_item_additional begin
//   // pragma uvmf custom class_item_additional end
  
//   // ****************************************************************************
//   covergroup data_mem_transaction_cg;
//     // pragma uvmf custom covergroup begin
//     // UVMF_CHANGE_ME : Add coverage bins, crosses, exclusions, etc. according to coverage needs.
//     option.auto_bin_max=1024;
//     option.per_instance=1;
//     complete_data: coverpoint coverage_trans.complete_data;
//     Data_dout: coverpoint coverage_trans.Data_dout;
//     Data_din: coverpoint coverage_trans.Data_din;
//     Data_rd: coverpoint coverage_trans.Data_rd;
//     Data_addr: coverpoint coverage_trans.Data_addr;
//     // pragma uvmf custom covergroup end
//   endgroup

//   // ****************************************************************************
//   // FUNCTION : new()
//   // This function is the standard SystemVerilog constructor.
//   //
//   function new(string name="", uvm_component parent=null);
//     super.new(name,parent);
//     data_mem_transaction_cg=new;
//     `uvm_warning("COVERAGE_MODEL_REVIEW", "A covergroup has been constructed which may need review because of either generation or re-generation with merging.  Please note that transaction variables added as a result of re-generation and merging are not automatically added to the covergroup.  Remove this warning after the covergroup has been reviewed.")
//   endfunction

//   // ****************************************************************************
//   // FUNCTION : build_phase()
//   // This function is the standard UVM build_phase.
//   //
//   function void build_phase(uvm_phase phase);
//     data_mem_transaction_cg.set_inst_name($sformatf("data_mem_transaction_cg_%s",get_full_name()));
//   endfunction

//   // ****************************************************************************
//   // FUNCTION: write (T t)
//   // This function is automatically executed when a transaction arrives on the
//   // analysis_export.  It copies values from the variables in the transaction 
//   // to local variables used to collect functional coverage.  
//   //
//   virtual function void write (T t);
//     `uvm_info("COV","Received transaction",UVM_HIGH);
//     coverage_trans = t;
//     data_mem_transaction_cg.sample();
//   endfunction

// endclass

// // pragma uvmf custom external begin
// // pragma uvmf custom external end

